`timescale 1ns / 1ps
module front_show(
//  HDMI IN PORT
//    input             pixclk_in,                            
    input             vs_in, 
    input             hs_in, 
    input             de_in,
//    input     [7:0]   r_in, 
//    input     [7:0]   g_in, 
//    input     [7:0]   b_in,
    input     [3:0]   led , 
//       
//    input      [10:0]  pixel_x,
//    input      [10:0]  pixel_y,
    input      [23:0]  front_colour,//������ɫ
    input      [23:0]  back_colour,//���ֱ�����ɫ
    input      [23:0]  default_colour,//Ĭ����ɫ
    input              pixel_clk,
    output             front_de,
    output reg [23:0]  pixel_data_out
    );
    parameter               H_TOTAL = 12'd1920;
    parameter               V_TOTAL = 12'd1080;
parameter front_xstart=16'd10;//�ַ�����ʼx����
parameter front_ystart=16'd10;//�ַ�����ʼy����  
parameter front_num=16'd5;//��ʾ����������
parameter front_width=8'd24;
parameter front_high=8'd24;
parameter front_len=1600;//24x24��ģӢ�ĳ����Ϊ24:12�������ַ����Ϊ4�����ص㣬���ʵ�ʳ���ΪW=12+4=16,H=24,W*H=16*24=384   
/*�ֿ�*/
reg [front_len-1:0]string_0 [front_num-1:0];
reg [front_len-1:0]used_string;
reg [11:0]        h_count = 'd0;
reg [11:0]        v_count = 'd0;
initial begin
string_0[0]=1600'h000000000000000000000000000000000000000000000000000000000000000006000000000E00000000FE0000007FFE000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000003E000000007F0000007FFFFF000000000000000000000000000000000000000000000000000000000000000000000000;/*"1"0*//*"0",0*/
string_0[1]=1600'h00000000000000000000000000000000000000000000000000000000000000007F0000001F87F8000078003E0001E0001F8003C0000FC007C00007C007E00007C007F00007C003F00007C00000000FC00000000F800000001F000000003C00000000F800000001E000000007800000001E000000007800000001E000000007800000001E000000003800006000E00000C003C00001C007000007C00FFFFFFFC00FFFFFFF800000000000000000000000000000000000000000000000000000000000000000000000;/*"2"0*/
string_0[2]=1600'h0000000000000000000000000000000000000000000000000000000000000000FC0000001F0FE00000F000F80001E0003E0003E0001F0003F0001F8003F0001F8001E0001F800000001F000000001F000000007C00000001F00000007F80000001FFC000000000F8000000001F000000000F8000000007C000000007E000000007E001C00007E007F00007E007F00007C007E0000F8003E0001F0001F0007C00003F07F0000001FE0000000000000000000000000000000000000000000000000000000000000000;/*"3"0*/
string_0[3]=1600'h0000000000000000000000000000000000000000000000000000000000000000007800000000F800000001F800000003F80000000EF80000001CF800000038F800000060F8000001C0F800000380F800000700F800000C00F800003800F800007000F80000C000F800018000F800070000F8000E0000F8001FFFFFFFF8000000F800000000F800000000F800000000F800000000F800000000F800000001F8000000FFFFF00000000000000000000000000000000000000000000000000000000000000000000000;/*"4"0*/
string_0[4]=1600'h00000000000000000000000000008000000003C007FFFFFFE0000038000000003800000000380000000030000000003000000000300000000030000000003000000000300000000030006000003000F03FFFFFFFF8000076000000007600000000660000000066000000006600000000E600000000C600000001C6000000018600000001860010000306001000070600100006060010000C0600100018060010003006001800E007003C018007FFFC070003FFF00C00000000300000000000000000000000000000;/*"��"0*/

//string[1]=384'h0000000000000000000002003E0006000600060006000600060006000600060006000600060006003FC0000000000000;/*"1",1*/
//string[2]=384'h000000000000000000001F00218040C060C060C000C00080018003000600040008001040204060407FC0000000000000;/*"2",2*/
//string[3]=384'h000000000000000000001E006300618061800180018003000E000180008000C000C060C060C061801F00000000000000;/*"3",3*/
//string[4]=384'h0000000000000000000001800180038005800580098011801180218041807FF0018001800180018007E0000000000000;/*"4",4*/
//string[5]=384'h000000000000000000003FC0200020002000200020002F00318020C000C000C060C060C0418021801F00000000000000;/*"5",5*/
//string[6]=384'h00000000000000000000078018C030C0300020006000678068C070606060606060602060304018C00F00000000000000;/*"6",6*/
//string[7]=384'h000000000000000000001FE0306020402080008000800100010002000200020006000600060006000600000000000000;/*"7",7*/
//string[8]=384'h000000000000000000001F8030C0606060606060304038C00F00138030C0606060606060606030C00F80000000000000;/*"8",8*/
//string[9]=384'h000000000000000000000F00308030C0604060606060606060E031601E60006000C000C0308031801E00000000000000;/*"9",9*/
//string[10]=384'h00000000000000000000FFC060C0602060206000610061007F006100610061006000600060006000F800000000000000;/*"F"10*/
//string[11]=384'h00000000000000000000FF0060C06060606060606060606061C07F00600060006000600060006000F800000000000000;/*"P"11*/
//string[12]=384'h000000000000000000000F001880304030402040600060006000600063F060C060C030C030C018C00F00000000000000;/*"G"12*/
//string[13]=384'h00000000000000000000060006000A000B00090009001100118010801F8020C020C0204040404060F0F0000000000000;/*"A"13*/
//string[14]=384'h000000000000000000000000040004000C000C007F800C000C000C000C000C000C000C000C400C400780000000000000;/*"t"14*/
//string[15]=384'h0000000000000000000000000000000000000000078018C01040306030603FE030003000182018400780000000000000;/*"e"15*/
//string[16]=384'h00000000000000000000000000000000000000000FC038C0304030401C000F0003C020C020C031C03F80000000000000;/*"s"16*/
//string[17]=384'h000000000000000000000000040004000C000C007F800C000C000C000C000C000C000C000C400C400780000000000000;/*"t"17*/
end
/*�ֿ�*/
reg [11:0]string_width = front_width;//�4095
wire [10:0]x_cnt;
wire [10:0]y_cnt;
assign front_de = (h_count >= front_xstart) && (h_count<(front_xstart+string_width)) && (v_count>=front_ystart) && (v_count<front_ystart+front_high) ;
assign x_cnt = h_count-front_xstart; //���ص�������ַ�������ʼ��ˮƽ����
assign y_cnt = v_count-front_ystart; //���ص�������ַ�������ʼ�㴹ֱ����/����ʱ��

always@(*)begin
case(led) 
4'b0001:used_string<=string_0[0];
4'b0010:used_string<=string_0[1];
4'b0100:used_string<=string_0[2];
4'b1000:used_string<=string_0[3];
default: used_string<=string_0[4];
endcase
end


always @(posedge pixel_clk ) 
begin    
        if(front_de)
        begin 
//            if(string[x_cnt/front_width][front_len-(x_cnt%front_width+(y_cnt-1)*front_width)]!=0)
              if(used_string[front_len-(x_cnt%front_width+(y_cnt-1)*front_width)]!=0)
                pixel_data_out <= front_colour;
            else
                pixel_data_out <= back_colour;
        end
        else
                pixel_data_out <= default_colour;                         
end    


   /* horizontal counter */
    always @(posedge pixel_clk)
    begin
        if (vs_in)
//        if (!rst_n|vs_in)
            h_count <= 'd0;
        else
        begin
            if ( (h_count < H_TOTAL - 1)&de_in   )
                h_count <= h_count + 1;
            else
                h_count <= 'd0;
        end
    end
    
    /* vertical counter */
    always @(posedge pixel_clk)
    begin
        if (vs_in)
//        if (!rst_n|vs_in)
            v_count <=  'd0;
        else
//        if (vs_in)
//            v_count <=  'd0;
//        else
        if (h_count == H_TOTAL - 1)
        begin
            if (v_count == V_TOTAL - 1)
                v_count <= 'd0;
            else
                v_count <= v_count + 1;
        end
    end


endmodule